// squares.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module squares (
		input  wire        clk_clk,              //      clk.clk
		output wire [41:0] hex_new_signal,       //      hex.new_signal
		input  wire [3:0]  keys_new_signal,      //     keys.new_signal
		output wire [9:0]  ledr_new_signal,      //     ledr.new_signal
		input  wire        ps2_conduit_end_clk,  //      ps2.conduit_end_clk
		input  wire        ps2_conduit_end_data, //         .conduit_end_data
		input  wire        reset_reset_n,        //    reset.reset_n
		input  wire [9:0]  switches_new_signal,  // switches.new_signal
		output wire        vga_CLK,              //      vga.CLK
		output wire        vga_HS,               //         .HS
		output wire        vga_VS,               //         .VS
		output wire        vga_BLANK,            //         .BLANK
		output wire        vga_SYNC,             //         .SYNC
		output wire [7:0]  vga_R,                //         .R
		output wire [7:0]  vga_G,                //         .G
		output wire [7:0]  vga_B                 //         .B
	);

	wire         game_0_avalon_streaming_source_valid;         // game_0:avalon_streaming_source_valid -> video_vga_controller_0:valid
	wire  [29:0] game_0_avalon_streaming_source_data;          // game_0:avalon_streaming_source_data -> video_vga_controller_0:data
	wire         game_0_avalon_streaming_source_ready;         // video_vga_controller_0:ready -> game_0:avalon_streaming_source_ready
	wire         game_0_avalon_streaming_source_startofpacket; // game_0:avalon_streaming_source_startofpacket -> video_vga_controller_0:startofpacket
	wire         game_0_avalon_streaming_source_endofpacket;   // game_0:avalon_streaming_source_endofpacket -> video_vga_controller_0:endofpacket
	wire         pll_0_outclk0_clk;                            // pll_0:outclk_0 -> game_0:clock_ps
	wire         video_pll_0_vga_clk_clk;                      // video_pll_0:vga_clk_clk -> [game_0:clock_vga, rst_controller:clk, video_vga_controller_0:clk]
	wire         rst_controller_reset_out_reset;               // rst_controller:reset_out -> [game_0:reset_reset, video_vga_controller_0:reset]

	game game_0 (
		.reset_reset                           (rst_controller_reset_out_reset),               //                   reset.reset
		.conduit_end_clk                       (ps2_conduit_end_clk),                          //             conduit_end.conduit_end_clk
		.conduit_end_data                      (ps2_conduit_end_data),                         //                        .conduit_end_data
		.avalon_streaming_source_data          (game_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.avalon_streaming_source_startofpacket (game_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.avalon_streaming_source_endofpacket   (game_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.avalon_streaming_source_valid         (game_0_avalon_streaming_source_valid),         //                        .valid
		.avalon_streaming_source_ready         (game_0_avalon_streaming_source_ready),         //                        .ready
		.clock_vga                             (video_pll_0_vga_clk_clk),                      //               clock_vga.clk
		.clock                                 (clk_clk),                                      //                clock_50.clk
		.clock_ps                              (pll_0_outclk0_clk),                            //                clock_ps.clk
		.conduit_end_1_new_signal              (ledr_new_signal),                              //           conduit_end_1.new_signal
		.conduit_end_2_new_signal              (hex_new_signal),                               //           conduit_end_2.new_signal
		.keys                                  (keys_new_signal),                              //                    keys.new_signal
		.switches                              (switches_new_signal)                           //                switches.new_signal
	);

	squares_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	squares_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                 //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),          //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk), //      vga_clk.clk
		.reset_source_reset ()                         // reset_source.reset
	);

	squares_video_vga_controller_0 video_vga_controller_0 (
		.clk           (video_pll_0_vga_clk_clk),                      //                clk.clk
		.reset         (rst_controller_reset_out_reset),               //              reset.reset
		.data          (game_0_avalon_streaming_source_data),          //    avalon_vga_sink.data
		.startofpacket (game_0_avalon_streaming_source_startofpacket), //                   .startofpacket
		.endofpacket   (game_0_avalon_streaming_source_endofpacket),   //                   .endofpacket
		.valid         (game_0_avalon_streaming_source_valid),         //                   .valid
		.ready         (game_0_avalon_streaming_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                      // external_interface.export
		.VGA_HS        (vga_HS),                                       //                   .export
		.VGA_VS        (vga_VS),                                       //                   .export
		.VGA_BLANK     (vga_BLANK),                                    //                   .export
		.VGA_SYNC      (vga_SYNC),                                     //                   .export
		.VGA_R         (vga_R),                                        //                   .export
		.VGA_G         (vga_G),                                        //                   .export
		.VGA_B         (vga_B)                                         //                   .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
