module dummy_entities();


endmodule