module game_logic();
	

endmodule