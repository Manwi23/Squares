module game_logic(
	output reg [6:0] address_write_om,
	output reg [10:0] data_write_om,
	output reg [6:0] address_read_om,
	input [10:0] data_read_om,
	input next_screen,
	output reg new_state,
	input clk
);
	

endmodule