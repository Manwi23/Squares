module operational_memory(
	input [6:0] address_write,
	input [10:0] data_write,
	input wren,
	input [6:0] address_read,
	output [10:0] data_read,
	input next_screen,
	input new_state,
	input clk
);



endmodule